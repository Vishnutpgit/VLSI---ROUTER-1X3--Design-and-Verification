package router_pkg ;
 
   import uvm_pkg::*;
   `include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "write_xtn.sv"
`include "router_src_agt_config.sv"    
`include "router_dst_agt_config.sv"
`include "router_env_config.sv"
`include "router_src_driver.sv"
`include "router_src_monitor.sv"
`include "router_src_sequencer.sv"
`include "router_src_agt.sv"
`include "router_src_agt_top.sv"
`include "router_src_sequence.sv"

`include "read_xtn.sv"
`include "router_dst_driver.sv"
`include "router_dst_monitor.sv"
`include "router_dst_sequencer.sv"
`include "router_dst_agt.sv"
`include "router_dst_agt_top.sv"
`include "router_dst_sequence.sv"


`include "router_v_sequencer.sv"
//`include "router_v_sequence.sv"
`include "router_sb.sv"

`include "router_env.sv"
`include "router_test.sv"


endpackage 
