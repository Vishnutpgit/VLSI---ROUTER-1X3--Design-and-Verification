class router_v_sequencer extends uvm_sequencer #(uvm_sequence_item) ;

 `uvm_component_utils(router_v_sequencer)

  router_src_sequencer src_seqrh[] ;
  router_dst_sequencer dst_seqrh[] ; 

extern function new(string name = "router_v_sequencer" , uvm_component parent = null);

endclass



function router_v_sequencer::new(string name = "router_v_sequencer" , uvm_component parent = null);
super.new(name,parent);
endfunction



